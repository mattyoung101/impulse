module multiplier(input logic [8:0] a, b, output logic[17:0] y);
    assign y = a * b;
endmodule