// This file is part of Impulse, the retro FPGA synthesizer
// Copyright (c) 2022 Matt Young. All rights reserved.

// Noise oscillator for Impulse
// This oscillator is based on a 16-bit maximal-period LFSR, sourced from:
// https://en.wikipedia.org/wiki/Linear-feedback_shift_register#Example_polynomials_for_maximal_LFSRs